`timescale 1ns/10ps
`define CYCLE_TIME 10



module PATTERN(
	clk,
	opA,
	opB,
	opM,
	out_data
);

//---------------------------------------------------------------------
// Input Output Declare
//---------------------------------------------------------------------
output reg	clk;
output reg [255:0]	opA,opB,opM;
input [255:0]	out_data;

//---------------------------------------------------------------------
// Register, parameter declaration
//---------------------------------------------------------------------
integer patcount;
parameter PATNUM = 10;

integer in_read,out_read;
integer i,j,a,gap;

integer counter;
integer curr_cycle, cycles, total_cycles;


//================================================================
// clock
//================================================================
always	#(`CYCLE_TIME/2.0) clk = ~clk;
initial	clk = 0;

reg [255:0]golden = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000101111101110011101011111001000011110100001100001000101;

initial begin
	opA = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011110111101111111110011000101100100001001101111101100101011;
	opB = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001110001101110101010011001100100010100110001110100011010;
	opM = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111010010010111101000110011010000001101100100000101000001;
	@(negedge clk);
	if(out_data!=golden) $display("Error!\n");
	else $display("Pass!!\n");
	$finish;
end


endmodule